`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:37:32 12/28/2014 
// Design Name: 
// Module Name:    bridge_sm 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bridge_sm(
    input GPS_I0,
    input GPS_I1,
    input GPS_Q0,
    input GPS_Q1,
    input MCU_CLK_25_000,
    output MCU_SCK,
    output MCU_SS,
    output MCU_MOSI
    );


endmodule
