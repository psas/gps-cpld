`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:43:04 12/28/2014 
// Design Name: 
// Module Name:    asynch_edge_detect 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module asynch_edge_detect(
    input SYNC_CLK_IN,
    input ASYNC_IN,
    output SYNC_OUT
    );


endmodule
